package dlx_types is
  subtype dlx_word is bit_vector(31 downto 0); 
  subtype half_word is bit_vector(15 downto 0);
  subtype byte is bit_vector(7 downto 0); 

  subtype alu_operation_code is bit_vector(3 downto 0); 
  subtype error_code is bit_vector(3 downto 0); 
  subtype register_index is bit_vector(4 downto 0); 

  subtype opcode_type is bit_vector(5 downto 0);
  subtype threeway_muxcode is bit_vector (1 downto 0);
  subtype func_code is bit_vector (5 downto 0);
end package dlx_types; 
